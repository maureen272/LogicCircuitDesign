// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sat Oct 07 11:56:02 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module control_unit (
    reset,clock,star,chk,sharp,count,
    ce,rw);

    input reset;
    input clock;
    input star;
    input chk;
    input sharp;
    input [1:0] count;
    tri0 reset;
    tri0 star;
    tri0 chk;
    tri0 sharp;
    tri0 [1:0] count;
    output ce;
    output rw;
    reg ce;
    reg rw;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or star or chk or sharp or count)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            ce <= 1'b0;
            rw <= 1'b0;
        end
        else begin
            ce <= 1'b0;
            rw <= 1'b0;
            case (fstate)
                state1: begin
                    if ((star == 1'b0))
                        reg_fstate <= state1;
                    else if ((star == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    rw <= 1'b0;

                    ce <= 1'b0;
                end
                state2: begin
                    if ((chk == 1'b0))
                        reg_fstate <= state2;
                    else if ((chk == 1'b1))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    rw <= 1'b0;

                    ce <= 1'b0;
                end
                state3: begin
                    if ((count[1:0] == 2'b11))
                        reg_fstate <= state4;
                    else if ((count[1:0] != 2'b11))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    rw <= 1'b1;

                    ce <= 1'b1;
                end
                state4: begin
                    if ((sharp == 1'b0))
                        reg_fstate <= state4;
                    else if ((sharp == 1'b1))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    rw <= 1'b0;

                    ce <= 1'b0;
                end
                state5: begin
                    if ((count[1:0] != 2'b11))
                        reg_fstate <= state5;
                    else if ((count[1:0] == 2'b11))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    rw <= 1'b0;

                    ce <= 1'b1;
                end
                default: begin
                    ce <= 1'bx;
                    rw <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // control_unit
